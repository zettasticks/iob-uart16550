//add primary io to system instance


   //UART16550
   output                   uart_txd,
   input                    uart_rxd,
   output                   uart_rts,
   input                    uart_cts,
